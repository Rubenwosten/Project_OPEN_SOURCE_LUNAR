* Analog block group 1 simulation
.subckt RL VinL Vout
*.ipin VinL
*.opin Vout
R1 Vout GND 1k m=1
R2 VinL Vout 1k m=1
.ends RL


Vnet7 net7 0 PWL(0n 0 0n -0.35714285714285715 0n -0.5 0n -0.35714285714285715 0n -0.5 0n -0.35714285714285715 0n -0.5 0n -0.35714285714285715 1n -0.5 1n -0.35714285714285715 1n 0.0714285714285714 2n -0.2142857142857143 2n 0.0714285714285714 3n 0.3571428571428571 4n 0.3571428571428571 5n 0.3571428571428571 6n 0.0714285714285714 7n -0.5 8n -0.5 9n -0.5 10n -0.5 11n -0.5 12n -0.2142857142857143 13n 0.3571428571428571 14n 0.3571428571428571 15n 0.3571428571428571 16n 0.0714285714285714 17n -0.5 18n -0.5 19n -0.5 20n -0.5 21n -0.5 22n -0.2142857142857143 23n 0.3571428571428571 24n 0.3571428571428571 25n 0.3571428571428571 26n 0.0714285714285714 27n -0.5 28n -0.5 29n -0.5 30n -0.5 31n -0.5 32n -0.2142857142857143 33n 0.3571428571428571 34n 0.3571428571428571 35n 0.3571428571428571 36n 0.0714285714285714 37n -0.5 38n -0.5 39n -0.5 40n -0.5 41n -0.5 42n -0.2142857142857143 43n 0.3571428571428571 44n 0.3571428571428571 45n 0.3571428571428571 46n 0.0714285714285714 47n -0.5 48n -0.5 49n -0.5)

X7 net7 VOUT RL

.control
   tran 50.0000p 50.0000n
   .probe
   wrdata VOUT.txt V(VOUT)
.endc
.end