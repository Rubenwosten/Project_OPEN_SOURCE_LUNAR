// inverter.v
module inverter (
    input wire a,
    output wire y
);
    assign y = ~a;
endmodule
