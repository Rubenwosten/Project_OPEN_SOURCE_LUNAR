* Analog block group 1 simulation
.subckt RL VinL Vout
*.ipin VinL
*.opin Vout
R1 Vout GND 1k m=1
R2 VinL Vout 1k m=1
.ends RL


Vnet7 net7 0 PWL(0n 0 0.0n -0.35714285714285715 0.01n -0.5 0.02n -0.35714285714285715 0.04n -0.5 0.08n -0.35714285714285715 0.16n -0.5 0.32n -0.35714285714285715 0.64n -0.5 0.98n -0.35714285714285715 1.37n 0.0714285714285714 1.73n -0.07142857142857145 2.38n 0.2142857142857143 3.17n 0.5 4.17n 0.5 5.17n 0.5 6.17n 0.2142857142857143 7.17n -0.35714285714285715 8.17n -0.35714285714285715 9.17n -0.35714285714285715 10.17n -0.35714285714285715 11.17n -0.35714285714285715 12.17n -0.07142857142857145 13.17n 0.5 14.17n 0.5 15.17n 0.5 16.17n 0.2142857142857143 17.17n -0.35714285714285715 18.17n -0.35714285714285715 19.17n -0.35714285714285715 20.17n -0.35714285714285715 21.17n -0.35714285714285715 22.17n -0.07142857142857145 23.17n 0.5 24.17n 0.5 25.17n 0.5 26.17n 0.2142857142857143 27.17n -0.35714285714285715 28.17n -0.35714285714285715 29.17n -0.35714285714285715 30.17n -0.35714285714285715 31.17n -0.35714285714285715 32.17n -0.07142857142857145 33.17n 0.5 34.17n 0.5 35.17n 0.5 36.17n 0.2142857142857143 37.17n -0.35714285714285715 38.17n -0.35714285714285715 39.17n -0.35714285714285715 40.17n -0.35714285714285715 41.17n -0.35714285714285715 42.17n -0.07142857142857145 43.17n 0.5 44.17n 0.5 45.17n 0.5 46.17n 0.2142857142857143 47.17n -0.35714285714285715 48.17n -0.35714285714285715 49.17n -0.35714285714285715 49.17n -0.35714285714285715)

X7 net7 VOUT RL

.control
   tran 50.0000p 50.0000n
   .probe
   wrdata VOUT.txt V(VOUT)
.endc
.end