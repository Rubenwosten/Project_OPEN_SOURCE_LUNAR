* Flattened netlist for RL

.subckt RL VINL VOUT
R1 VOUT GND 1k
R2 VINL VOUT 1k
.ends RL
